--------------------------------------------------------------------------------
-- Title       : Testbed for FSK receiver on Altera DE1-SoC
-- Project     : FPGA Based Digital Signal Processing
--               FH OÖ Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: TbdRxFskBasic-e.vhd 733 2017-12-04 02:28:35Z mroland $
-- Authors     : Markus Pfaff, Linz/Austria, Copyright (c) 2003-2005
--               Michael Roland, Hagenberg/Austria, Copyright (c) 2011-2017
--------------------------------------------------------------------------------
-- Description : Decoded output to LED
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- fixed_pkg resides in the library ieee since VHDL-2008 (QuestaSim backports
-- this to VHDL-93 too). However, Quartus (as of version 13.0sp1) still does
-- not have native support for ieee.fixed_pkg. Therefore, we provide the
-- VHDL-93 compatibility versions as part of this excercise. These must be
-- compiled into the are located in the library ieee_proposed. Include them in
-- your Config.tcl and don't forget to set the ExtraLibraries and TargetLibrary
-- parameters to compile them into the right library (ieee_proposed) with fhlow.
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
-- In future (when both QuestaSim and Quartus support the VHDL-2008
-- ieee.fixed_pkg) simply use:
--use ieee.fixed_float_types.all;
--use ieee.fixed_pkg.all;

use work.Global.all;
use work.DefinitionsCodec.all;
use work.ParamCodec.all;
use work.DefinitionsFsk.all;

entity TbdRxFskBasic is

  generic (
    gClkFrequency      : natural            := cDefaultClkFrequency;
    gAudioBitWidth     : natural            := cDefaultAudioBitWidth;
    gSampleRate        : natural            := cDefaultSampleRate;
    -- Rx parameters
    gCoefWidth         : natural            := cFskFilterCoefWidth;
    -- The values used as filter coefficients. The number of those
    -- coefficients determines the number of taps the filter has.
    gChannelBandpasses : aSetOfRxBandpasses := (
      0               => (Bandpass0 => (-0.003244924172431670000000, 0.002951979629087140000000, 0.002163282781621110000000, 0.001284449151587530000000, 0.000473218108479618000000, 0.000202807760776979000000, 0.000383081325912072000000, 0.000518286499763391000000, 0.000247876152060752000000, -0.000135205173851319000000, -0.000180273565135093000000, 0.000090136782567546300000, 0.000247876152060752000000, 0.000090136782567546300000, -0.000112670978209433000000, -0.000112670978209433000000, 0.000022534195641886600000, 0.000045068391283773100000, 0.000000000000000000000000, 0.000022534195641886600000, 0.000090136782567546300000, -0.000022534195641886600000, -0.000202807760776979000000, -0.000135205173851319000000, 0.000247876152060752000000, 0.000360547130270185000000, -0.000067602586925659700000, -0.000563354891047164000000, -0.000315478738986412000000, 0.000518286499763391000000, 0.000766162651824143000000, -0.000112670978209433000000, -0.001014038803884900000000, -0.000563354891047164000000, 0.000833765238749803000000, 0.001261914955945650000000, -0.000135205173851319000000, -0.001577393694932060000000, -0.000901367825675463000000, 0.001216846564661870000000, 0.001847804042634700000000, -0.000157739369493206000000, -0.002230885368546770000000, -0.001306983347229420000000, 0.001644996281857720000000, 0.002568898303175070000000, -0.000135205173851319000000, -0.002951979629087140000000, -0.001802735651350930000000, 0.002095680194695450000000, 0.003380129346282980000000, -0.000090136782567546300000, -0.003785744867836940000000, -0.002388624738039980000000, 0.002568898303175070000000, 0.004281497171958450000000, 0.000000000000000000000000, -0.004642044302228630000000, -0.003042116411654690000000, 0.003042116411654690000000, 0.005273001780201460000000, 0.000135205173851319000000, -0.005565946323545980000000, -0.003763210672195060000000, 0.003515334520134300000000, 0.006309574779728240000000, 0.000338012934628298000000, -0.006512382540505220000000, -0.004574441715302970000000, 0.003966018432972040000000, 0.007413750366180680000000, 0.000585889086689051000000, -0.007458818757464450000000, -0.005408206954052780000000, 0.004371633954525990000000, 0.008517925952633120000000, 0.000878833630033576000000, -0.008360186583139920000000, -0.006287040584086350000000, 0.004732181084796180000000, 0.009599567343443680000000, 0.001216846564661870000000, -0.009239020213173490000000, -0.007188408409761810000000, 0.005002591432498820000000, 0.010658674538612300000000, 0.001622462086215830000000, -0.010005182864997600000000, -0.008067242039795390000000, 0.005205399193275800000000, 0.011650179146855400000000, 0.002050611803411680000000, -0.010703742929896100000000, -0.008901007278545190000000, 0.005340604367127120000000, 0.012529012776888900000000, 0.002501295716249410000000, -0.011267097820943300000000, -0.009712238321653110000000, 0.005363138562769000000000, 0.013317709624355000000000, 0.002951979629087140000000, -0.011695247538139100000000, -0.010410798386551600000000, 0.005295535975843340000000, 0.013926132906685900000000, 0.003425197737566760000000, -0.011965657885841800000000, -0.011019221668882500000000, 0.005160330801992020000000, 0.014399351015165500000000, 0.003853347454762600000000, -0.012078328864051200000000, -0.011514973973004000000000, 0.004934988845573160000000, 0.014669761362868200000000, 0.004258962976316560000000, -0.012055794668409300000000, -0.011852986907632300000000, 0.004642044302228630000000, 0.014759898145435700000000, 0.004642044302228630000000, -0.011852986907632300000000, -0.012055794668409300000000, 0.004258962976316560000000, 0.014669761362868200000000, 0.004934988845573160000000, -0.011514973973004000000000, -0.012078328864051200000000, 0.003853347454762600000000, 0.014399351015165500000000, 0.005160330801992020000000, -0.011019221668882500000000, -0.011965657885841800000000, 0.003425197737566760000000, 0.013926132906685900000000, 0.005295535975843340000000, -0.010410798386551600000000, -0.011695247538139100000000, 0.002951979629087140000000, 0.013317709624355000000000, 0.005363138562769000000000, -0.009712238321653110000000, -0.011267097820943300000000, 0.002501295716249410000000, 0.012529012776888900000000, 0.005340604367127120000000, -0.008901007278545190000000, -0.010703742929896100000000, 0.002050611803411680000000, 0.011650179146855400000000, 0.005205399193275800000000, -0.008067242039795390000000, -0.010005182864997600000000, 0.001622462086215830000000, 0.010658674538612300000000, 0.005002591432498820000000, -0.007188408409761810000000, -0.009239020213173490000000, 0.001216846564661870000000, 0.009599567343443680000000, 0.004732181084796180000000, -0.006287040584086350000000, -0.008360186583139920000000, 0.000878833630033576000000, 0.008517925952633120000000, 0.004371633954525990000000, -0.005408206954052780000000, -0.007458818757464450000000, 0.000585889086689051000000, 0.007413750366180680000000, 0.003966018432972040000000, -0.004574441715302970000000, -0.006512382540505220000000, 0.000338012934628298000000, 0.006309574779728240000000, 0.003515334520134300000000, -0.003763210672195060000000, -0.005565946323545980000000, 0.000135205173851319000000, 0.005273001780201460000000, 0.003042116411654690000000, -0.003042116411654690000000, -0.004642044302228630000000, 0.000000000000000000000000, 0.004281497171958450000000, 0.002568898303175070000000, -0.002388624738039980000000, -0.003785744867836940000000, -0.000090136782567546300000, 0.003380129346282980000000, 0.002095680194695450000000, -0.001802735651350930000000, -0.002951979629087140000000, -0.000135205173851319000000, 0.002568898303175070000000, 0.001644996281857720000000, -0.001306983347229420000000, -0.002230885368546770000000, -0.000157739369493206000000, 0.001847804042634700000000, 0.001216846564661870000000, -0.000901367825675463000000, -0.001577393694932060000000, -0.000135205173851319000000, 0.001261914955945650000000, 0.000833765238749803000000, -0.000563354891047164000000, -0.001014038803884900000000, -0.000112670978209433000000, 0.000766162651824143000000, 0.000518286499763391000000, -0.000315478738986412000000, -0.000563354891047164000000, -0.000067602586925659700000, 0.000360547130270185000000, 0.000247876152060752000000, -0.000135205173851319000000, -0.000202807760776979000000, -0.000022534195641886600000, 0.000090136782567546300000, 0.000022534195641886600000, 0.000000000000000000000000, 0.000045068391283773100000, 0.000022534195641886600000, -0.000112670978209433000000, -0.000112670978209433000000, 0.000090136782567546300000, 0.000247876152060752000000, 0.000090136782567546300000, -0.000180273565135093000000, -0.000135205173851319000000, 0.000247876152060752000000, 0.000518286499763391000000, 0.000383081325912072000000, 0.000202807760776979000000, 0.000473218108479618000000, 0.001284449151587530000000, 0.002163282781621110000000, 0.002951979629087140000000, -0.003244924172431670000000),
-- band pass for Channel 0/freq. 0 all u
            Bandpass1 => (-0.004418394950405770000000, -0.001127141568981060000000, 0.001330027051397660000000, -0.001172227231740310000000, 0.000676284941388638000000, -0.000338142470694319000000, 0.000450856627592426000000, -0.000743913435527502000000, 0.000743913435527502000000, -0.000383228133453562000000, 0.000067628494138863800000, -0.000135256988277728000000, 0.000360685302073941000000, -0.000428313796212804000000, 0.000225428313796213000000, -0.000045085662759242600000, 0.000067628494138863800000, -0.000135256988277728000000, 0.000135256988277728000000, -0.000090171325518485100000, 0.000135256988277728000000, -0.000202885482416592000000, 0.000067628494138863800000, 0.000180342651036970000000, -0.000180342651036970000000, -0.000202885482416592000000, 0.000518485121731289000000, -0.000202885482416592000000, -0.000473399458972047000000, 0.000631199278629396000000, 0.000135256988277728000000, -0.000924256086564473000000, 0.000586113615870153000000, 0.000653742110009017000000, -0.001194770063119930000000, 0.000157799819657349000000, 0.001307484220018030000000, -0.001217312894499550000000, -0.000586113615870153000000, 0.001848512173128950000000, -0.000766456266907124000000, -0.001555455365193870000000, 0.002073940486925160000000, 0.000180342651036970000000, -0.002479711451758340000000, 0.001690712353471600000000, 0.001487826871055000000000, -0.003020739404869250000000, 0.000631199278629396000000, 0.002885482416591520000000, -0.002885482416591520000000, -0.001014427412082960000000, 0.003922452660054100000000, -0.001848512173128950000000, -0.002908025247971150000000, 0.004215509467989180000000, 0.000000000000000000000000, -0.004576194770063120000000, 0.003426510369702430000000, 0.002389540126239860000000, -0.005477908025247970000000, 0.001532912533814250000000, 0.004756537421100090000000, -0.005184851217312890000000, -0.001239855725879170000000, 0.006469792605951310000000, -0.003471596032461680000000, -0.004305680793507660000000, 0.006898106402164110000000, -0.000541027953110911000000, -0.006898106402164110000000, 0.005680793507664560000000, 0.003088367899008120000000, -0.008295761947700630000000, 0.002862939585211900000000, 0.006605049594229040000000, -0.007889990982867450000000, -0.001127141568981060000000, 0.009084761045987380000000, -0.005522993688007210000000, -0.005455365193868350000000, 0.009761045987376010000000, -0.001510369702434630000000, -0.009062218214607750000000, 0.008205590622182150000000, 0.003403967538322810000000, -0.011023444544634800000000, 0.004553651938683500000000, 0.008070333633904420000000, -0.010617673579801600000000, -0.000586113615870153000000, 0.011361587015329100000000, -0.007709648331830480000000, -0.006064021641118120000000, 0.012353471596032500000000, -0.002772768259693420000000, -0.010640216411181200000000, 0.010595130748422000000000, 0.003178539224526600000000, -0.013142470694319200000000, 0.006311992786293960000000, 0.008836789900811540000000, -0.012849413886384100000000, 0.000338142470694319000000, 0.012826871055004500000000, -0.009648331830477910000000, -0.006018935978358880000000, 0.014134355275022500000000, -0.004147880973850320000000, -0.011316501352569900000000, 0.012376014427412100000000, 0.002479711451758340000000, -0.014269612263300300000000, 0.007822362488728590000000, 0.008724075743913440000000, -0.014156898106402200000000, 0.001442741208295760000000, 0.013187556357078400000000, -0.010955816050495900000000, -0.005320108205590620000000, 0.014788097385031600000000, -0.005320108205590620000000, -0.010955816050495900000000, 0.013187556357078400000000, 0.001442741208295760000000, -0.014156898106402200000000, 0.008724075743913440000000, 0.007822362488728590000000, -0.014269612263300300000000, 0.002479711451758340000000, 0.012376014427412100000000, -0.011316501352569900000000, -0.004147880973850320000000, 0.014134355275022500000000, -0.006018935978358880000000, -0.009648331830477910000000, 0.012826871055004500000000, 0.000338142470694319000000, -0.012849413886384100000000, 0.008836789900811540000000, 0.006311992786293960000000, -0.013142470694319200000000, 0.003178539224526600000000, 0.010595130748422000000000, -0.010640216411181200000000, -0.002772768259693420000000, 0.012353471596032500000000, -0.006064021641118120000000, -0.007709648331830480000000, 0.011361587015329100000000, -0.000586113615870153000000, -0.010617673579801600000000, 0.008070333633904420000000, 0.004553651938683500000000, -0.011023444544634800000000, 0.003403967538322810000000, 0.008205590622182150000000, -0.009062218214607750000000, -0.001510369702434630000000, 0.009761045987376010000000, -0.005455365193868350000000, -0.005522993688007210000000, 0.009084761045987380000000, -0.001127141568981060000000, -0.007889990982867450000000, 0.006605049594229040000000, 0.002862939585211900000000, -0.008295761947700630000000, 0.003088367899008120000000, 0.005680793507664560000000, -0.006898106402164110000000, -0.000541027953110911000000, 0.006898106402164110000000, -0.004305680793507660000000, -0.003471596032461680000000, 0.006469792605951310000000, -0.001239855725879170000000, -0.005184851217312890000000, 0.004756537421100090000000, 0.001532912533814250000000, -0.005477908025247970000000, 0.002389540126239860000000, 0.003426510369702430000000, -0.004576194770063120000000, 0.000000000000000000000000, 0.004215509467989180000000, -0.002908025247971150000000, -0.001848512173128950000000, 0.003922452660054100000000, -0.001014427412082960000000, -0.002885482416591520000000, 0.002885482416591520000000, 0.000631199278629396000000, -0.003020739404869250000000, 0.001487826871055000000000, 0.001690712353471600000000, -0.002479711451758340000000, 0.000180342651036970000000, 0.002073940486925160000000, -0.001555455365193870000000, -0.000766456266907124000000, 0.001848512173128950000000, -0.000586113615870153000000, -0.001217312894499550000000, 0.001307484220018030000000, 0.000157799819657349000000, -0.001194770063119930000000, 0.000653742110009017000000, 0.000586113615870153000000, -0.000924256086564473000000, 0.000135256988277728000000, 0.000631199278629396000000, -0.000473399458972047000000, -0.000202885482416592000000, 0.000518485121731289000000, -0.000202885482416592000000, -0.000180342651036970000000, 0.000180342651036970000000, 0.000067628494138863800000, -0.000202885482416592000000, 0.000135256988277728000000, -0.000090171325518485100000, 0.000135256988277728000000, -0.000135256988277728000000, 0.000067628494138863800000, -0.000045085662759242600000, 0.000225428313796213000000, -0.000428313796212804000000, 0.000360685302073941000000, -0.000135256988277728000000, 0.000067628494138863800000, -0.000383228133453562000000, 0.000743913435527502000000, -0.000743913435527502000000, 0.000450856627592426000000, -0.000338142470694319000000, 0.000676284941388638000000, -0.001172227231740310000000, 0.001330027051397660000000, -0.001127141568981060000000, -0.004418394950405770000000)),
-- band pass for Channel 0/freq. 1 all o
      1               => (Bandpass0 => (-0.000410162925828871000000, 0.005149823402073600000000, 0.000569670730317876000000, -0.000091147316850860200000, -0.000319015608978011000000, -0.000205081462914435000000, 0.000091147316850860200000, 0.000296228779765296000000, 0.000205081462914435000000, -0.000068360487638145200000, -0.000250655121339866000000, -0.000182294633701720000000, 0.000045573658425430100000, 0.000182294633701720000000, 0.000113934146063575000000, -0.000022786829212715100000, -0.000068360487638145200000, -0.000022786829212715100000, 0.000000000000000000000000, -0.000045573658425430100000, -0.000091147316850860200000, 0.000000000000000000000000, 0.000205081462914435000000, 0.000250655121339866000000, 0.000000000000000000000000, -0.000364589267403441000000, -0.000455736584254301000000, -0.000022786829212715100000, 0.000569670730317876000000, 0.000683604876381452000000, 0.000091147316850860200000, -0.000774752193232312000000, -0.000979833656146747000000, -0.000182294633701720000000, 0.000979833656146747000000, 0.001321636094337470000000, 0.000296228779765296000000, -0.001207701948273900000000, -0.001686225361740910000000, -0.000455736584254301000000, 0.001435570240401050000000, 0.002119175116782500000000, 0.000683604876381452000000, -0.001663438532528200000000, -0.002574911701036800000000, -0.000934259997721317000000, 0.001868519995442630000000, 0.003076221943716530000000, 0.001253275606699330000000, -0.002050814629144350000000, -0.003623105844821690000000, -0.001617864874102770000000, 0.002210322433633360000000, 0.004169989745926860000000, 0.002050814629144350000000, -0.002347043408909650000000, -0.004762447305457450000000, -0.002552124871824090000000, 0.002438190725760510000000, 0.005354904864988040000000, 0.003099008772929250000000, -0.002460977554973230000000, -0.005947362424518630000000, -0.003691466332459840000000, 0.002460977554973230000000, 0.006562606813261940000000, 0.004329497550415860000000, -0.002369830238122370000000, -0.007132277543579810000000, -0.005035889256010030000000, 0.002233109262846080000000, 0.007701948273897690000000, 0.005765067790816910000000, -0.002028027799931640000000, -0.008226045345790130000000, -0.006539819984049220000000, 0.001754585849379060000000, 0.008704568759257150000000, 0.007314572177281530000000, -0.001412783411188330000000, -0.009137518514298740000000, -0.008112111199726560000000, 0.001002620485359460000000, 0.009502107781702180000000, 0.008909650222171590000000, -0.000546883901105161000000, -0.009821123390680190000000, -0.009707189244616610000000, 0.000000000000000000000000, 0.010048991682807300000000, 0.010481941437848900000000, 0.000592457559530591000000, -0.010185712658083600000000, -0.011233906801868500000000, -0.001230488777486610000000, 0.010254073145721800000000, 0.011940298507462700000000, 0.001914093653868060000000, -0.010231286316509100000000, -0.012578329725418700000000, -0.002643272188674950000000, 0.010117352170445500000000, 0.013170787284949300000000, 0.003372450723481830000000, -0.009912270707531050000000, -0.013694884356841700000000, -0.004124416087501420000000, 0.009616041927765750000000, 0.014127834111883300000000, 0.004876381451521020000000, -0.009228665831149600000000, -0.014469636550074100000000, -0.005628346815540620000000, 0.008772929246895300000000, 0.014720291671413900000000, 0.006334738521134780000000, -0.008248832175002850000000, -0.014857012646690200000000, -0.007018343397516240000000, 0.007656374615472260000000, 0.014925373134328400000000, 0.007656374615472260000000, -0.007018343397516240000000, -0.014857012646690200000000, -0.008248832175002850000000, 0.006334738521134780000000, 0.014720291671413900000000, 0.008772929246895300000000, -0.005628346815540620000000, -0.014469636550074100000000, -0.009228665831149600000000, 0.004876381451521020000000, 0.014127834111883300000000, 0.009616041927765750000000, -0.004124416087501420000000, -0.013694884356841700000000, -0.009912270707531050000000, 0.003372450723481830000000, 0.013170787284949300000000, 0.010117352170445500000000, -0.002643272188674950000000, -0.012578329725418700000000, -0.010231286316509100000000, 0.001914093653868060000000, 0.011940298507462700000000, 0.010254073145721800000000, -0.001230488777486610000000, -0.011233906801868500000000, -0.010185712658083600000000, 0.000592457559530591000000, 0.010481941437848900000000, 0.010048991682807300000000, 0.000000000000000000000000, -0.009707189244616610000000, -0.009821123390680190000000, -0.000546883901105161000000, 0.008909650222171590000000, 0.009502107781702180000000, 0.001002620485359460000000, -0.008112111199726560000000, -0.009137518514298740000000, -0.001412783411188330000000, 0.007314572177281530000000, 0.008704568759257150000000, 0.001754585849379060000000, -0.006539819984049220000000, -0.008226045345790130000000, -0.002028027799931640000000, 0.005765067790816910000000, 0.007701948273897690000000, 0.002233109262846080000000, -0.005035889256010030000000, -0.007132277543579810000000, -0.002369830238122370000000, 0.004329497550415860000000, 0.006562606813261940000000, 0.002460977554973230000000, -0.003691466332459840000000, -0.005947362424518630000000, -0.002460977554973230000000, 0.003099008772929250000000, 0.005354904864988040000000, 0.002438190725760510000000, -0.002552124871824090000000, -0.004762447305457450000000, -0.002347043408909650000000, 0.002050814629144350000000, 0.004169989745926860000000, 0.002210322433633360000000, -0.001617864874102770000000, -0.003623105844821690000000, -0.002050814629144350000000, 0.001253275606699330000000, 0.003076221943716530000000, 0.001868519995442630000000, -0.000934259997721317000000, -0.002574911701036800000000, -0.001663438532528200000000, 0.000683604876381452000000, 0.002119175116782500000000, 0.001435570240401050000000, -0.000455736584254301000000, -0.001686225361740910000000, -0.001207701948273900000000, 0.000296228779765296000000, 0.001321636094337470000000, 0.000979833656146747000000, -0.000182294633701720000000, -0.000979833656146747000000, -0.000774752193232312000000, 0.000091147316850860200000, 0.000683604876381452000000, 0.000569670730317876000000, -0.000022786829212715100000, -0.000455736584254301000000, -0.000364589267403441000000, 0.000000000000000000000000, 0.000250655121339866000000, 0.000205081462914435000000, 0.000000000000000000000000, -0.000091147316850860200000, -0.000045573658425430100000, 0.000000000000000000000000, -0.000022786829212715100000, -0.000068360487638145200000, -0.000022786829212715100000, 0.000113934146063575000000, 0.000182294633701720000000, 0.000045573658425430100000, -0.000182294633701720000000, -0.000250655121339866000000, -0.000068360487638145200000, 0.000205081462914435000000, 0.000296228779765296000000, 0.000091147316850860200000, -0.000205081462914435000000, -0.000319015608978011000000, -0.000091147316850860200000, 0.000569670730317876000000, 0.005149823402073600000000, -0.000410162925828871000000),
-- band pass for Channel 1/freq. 0, own u
            Bandpass1 => (-0.000660486938301410000000, 0.005101692213086750000000, 0.000637711526635844000000, -0.000250529528321224000000, 0.000068326234996697600000, 0.000296080351652356000000, -0.000159427881658961000000, -0.000250529528321224000000, 0.000204978704990093000000, 0.000159427881658961000000, -0.000227754116655659000000, -0.000091101646662263400000, 0.000204978704990093000000, 0.000000000000000000000000, -0.000159427881658961000000, 0.000022775411665565900000, 0.000068326234996697600000, -0.000022775411665565900000, 0.000000000000000000000000, -0.000045550823331131700000, -0.000068326234996697600000, 0.000136652469993395000000, 0.000068326234996697600000, -0.000296080351652356000000, 0.000000000000000000000000, 0.000432732821645751000000, -0.000136652469993395000000, -0.000523834468308015000000, 0.000364406586649054000000, 0.000569385291639146000000, -0.000660486938301410000000, -0.000501059056642449000000, 0.000979342701619332000000, 0.000273304939986790000000, -0.001275423053271690000000, 0.000068326234996697600000, 0.001480401758261780000000, -0.000546609879973581000000, -0.001548727993258480000000, 0.001138770583278290000000, 0.001434850934930650000000, -0.001753706698248570000000, -0.001093219759947160000000, 0.002323091989887720000000, 0.000501059056642449000000, -0.002778600223199030000000, 0.000296080351652356000000, 0.003006354339854690000000, -0.001252647641606120000000, -0.002960803516523560000000, 0.002300316578222150000000, 0.002550846106543380000000, -0.003325210103172620000000, -0.001776482109914140000000, 0.004167900334798550000000, 0.000660486938301410000000, -0.004760061038103260000000, 0.000728813173298107000000, 0.004942264331427790000000, -0.002300316578222150000000, -0.004623408568109870000000, 0.003871819983146200000000, 0.003803493748149500000000, -0.005306670918076840000000, -0.002459744459881110000000, 0.006422666089689570000000, 0.000660486938301410000000, -0.007037602204659850000000, 0.001412075523265080000000, 0.007060377616325420000000, -0.003644065866490540000000, -0.006377115266358440000000, 0.005762179151388160000000, 0.004987815154758920000000, -0.007584212084633430000000, -0.002960803516523560000000, 0.008859635137905120000000, 0.000455508233311317000000, -0.009429020429544270000000, 0.002345867401553280000000, 0.009132940077891910000000, -0.005192793859749010000000, -0.007971394082948050000000, 0.007789190789623520000000, 0.005967157856378250000000, -0.009884528662855580000000, -0.003234108456510350000000, 0.011205502539458400000000, 0.000000000000000000000000, -0.011592684537773000000000, 0.003461862573166010000000, 0.010909422187806000000000, -0.006809848088004190000000, -0.009201266312888610000000, 0.009725100781196620000000, 0.006559318559682970000000, -0.011934315712756500000000, -0.003165782221513650000000, 0.013164187942697100000000, -0.000660486938301410000000, -0.013255289589359300000000, 0.004600633156444300000000, 0.012139294417746600000000, -0.008267474434600410000000, -0.009907304074521150000000, 0.011342155009451800000000, 0.006695971029676360000000, -0.013460268294349400000000, -0.002801375634864600000000, 0.014462386407634300000000, -0.001434850934930650000000, -0.014189081467647500000000, 0.005625526681394770000000, 0.012640353474389000000000, -0.009383469606213130000000, -0.009952854897852280000000, 0.012344273122736700000000, 0.006354339854692870000000, -0.014257407702644200000000, -0.002186439519894320000000, 0.014917894640945600000000, -0.002186439519894320000000, -0.014257407702644200000000, 0.006354339854692870000000, 0.012344273122736700000000, -0.009952854897852280000000, -0.009383469606213130000000, 0.012640353474389000000000, 0.005625526681394770000000, -0.014189081467647500000000, -0.001434850934930650000000, 0.014462386407634300000000, -0.002801375634864600000000, -0.013460268294349400000000, 0.006695971029676360000000, 0.011342155009451800000000, -0.009907304074521150000000, -0.008267474434600410000000, 0.012139294417746600000000, 0.004600633156444300000000, -0.013255289589359300000000, -0.000660486938301410000000, 0.013164187942697100000000, -0.003165782221513650000000, -0.011934315712756500000000, 0.006559318559682970000000, 0.009725100781196620000000, -0.009201266312888610000000, -0.006809848088004190000000, 0.010909422187806000000000, 0.003461862573166010000000, -0.011592684537773000000000, 0.000000000000000000000000, 0.011205502539458400000000, -0.003234108456510350000000, -0.009884528662855580000000, 0.005967157856378250000000, 0.007789190789623520000000, -0.007971394082948050000000, -0.005192793859749010000000, 0.009132940077891910000000, 0.002345867401553280000000, -0.009429020429544270000000, 0.000455508233311317000000, 0.008859635137905120000000, -0.002960803516523560000000, -0.007584212084633430000000, 0.004987815154758920000000, 0.005762179151388160000000, -0.006377115266358440000000, -0.003644065866490540000000, 0.007060377616325420000000, 0.001412075523265080000000, -0.007037602204659850000000, 0.000660486938301410000000, 0.006422666089689570000000, -0.002459744459881110000000, -0.005306670918076840000000, 0.003803493748149500000000, 0.003871819983146200000000, -0.004623408568109870000000, -0.002300316578222150000000, 0.004942264331427790000000, 0.000728813173298107000000, -0.004760061038103260000000, 0.000660486938301410000000, 0.004167900334798550000000, -0.001776482109914140000000, -0.003325210103172620000000, 0.002550846106543380000000, 0.002300316578222150000000, -0.002960803516523560000000, -0.001252647641606120000000, 0.003006354339854690000000, 0.000296080351652356000000, -0.002778600223199030000000, 0.000501059056642449000000, 0.002323091989887720000000, -0.001093219759947160000000, -0.001753706698248570000000, 0.001434850934930650000000, 0.001138770583278290000000, -0.001548727993258480000000, -0.000546609879973581000000, 0.001480401758261780000000, 0.000068326234996697600000, -0.001275423053271690000000, 0.000273304939986790000000, 0.000979342701619332000000, -0.000501059056642449000000, -0.000660486938301410000000, 0.000569385291639146000000, 0.000364406586649054000000, -0.000523834468308015000000, -0.000136652469993395000000, 0.000432732821645751000000, 0.000000000000000000000000, -0.000296080351652356000000, 0.000068326234996697600000, 0.000136652469993395000000, -0.000068326234996697600000, -0.000045550823331131700000, 0.000000000000000000000000, -0.000022775411665565900000, 0.000068326234996697600000, 0.000022775411665565900000, -0.000159427881658961000000, 0.000000000000000000000000, 0.000204978704990093000000, -0.000091101646662263400000, -0.000227754116655659000000, 0.000159427881658961000000, 0.000204978704990093000000, -0.000250529528321224000000, -0.000159427881658961000000, 0.000296080351652356000000, 0.000068326234996697600000, -0.000250529528321224000000, 0.000637711526635844000000, 0.005101692213086750000000, -0.000660486938301410000000)));
-- band pass for Channel 1/freq. 1 own o
    gLowpass           : aSetOfFactors      := (-0.004856389621201610000000, 0.002802830581379210000000, 0.003274594144581660000000, 0.004356875260163730000000, 0.005855418343277370000000, 0.007770223393922580000000, 0.010018038018593000000000, 0.012543360621617900000000, 0.015346191202997100000000, 0.018343277369224400000000, 0.021479117524628800000000, 0.024725960871375100000000, 0.027972804218121300000000, 0.031164145969196600000000, 0.034216733731094800000000, 0.037047315110309400000000, 0.039572637713334300000000, 0.041764950742333800000000, 0.043513251005966400000000, 0.044817538504232000000000, 0.045622311641459700000000, 0.045872068821978600000000, 0.045622311641459700000000, 0.044817538504232000000000, 0.043513251005966400000000, 0.041764950742333800000000, 0.039572637713334300000000, 0.037047315110309400000000, 0.034216733731094800000000, 0.031164145969196600000000, 0.027972804218121300000000, 0.024725960871375100000000, 0.021479117524628800000000, 0.018343277369224400000000, 0.015346191202997100000000, 0.012543360621617900000000, 0.010018038018593000000000, 0.007770223393922580000000, 0.005855418343277370000000, 0.004356875260163730000000, 0.003274594144581660000000, 0.002802830581379210000000, -0.004856389621201610000000)
-- low pass
    );

  port (
    iClk         : in std_ulogic;
    inResetAsync : in std_ulogic;

    -- User interface
    iSwitch  : in  std_ulogic_vector(9 downto 0);  -- active high
    inButton : in  std_ulogic_vector(3 downto 1);  -- active low
    oSEG0    : out std_ulogic_vector(6 downto 0);  -- active low
    oSEG1    : out std_ulogic_vector(6 downto 0);  -- active low
    oSEG2    : out std_ulogic_vector(6 downto 0);  -- active low
    oSEG3    : out std_ulogic_vector(6 downto 0);  -- active low
    oSEG4    : out std_ulogic_vector(6 downto 0);  -- active low
    oSEG5    : out std_ulogic_vector(6 downto 0);  -- active low
    oLed     : out std_ulogic_vector(9 downto 0);  -- active high

    -- Audio codec
    oI2cSclk  : out   std_ulogic;
    ioI2cSdin : inout std_logic;

    oMclk : out std_ulogic;

    oBclk   : out std_ulogic;
    iADCdat : in  std_ulogic;
    oDACdat : out std_ulogic;
    oADClrc : out std_ulogic;
    oDAClrc : out std_ulogic);

end TbdRxFskBasic;
