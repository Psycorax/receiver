--------------------------------------------------------------------------------
-- Title       : Testbench for design "DspFir"
-- Project     : FPGA Based Digital Signal Processing
--               FH OÖ Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: tbDspFir-Bhv-ea.vhd 711 2017-11-03 18:22:43Z mroland $
-- Authors     : Markus Pfaff, Linz/Austria, Copyright (c) 2003-2005
--               Michael Roland, Hagenberg/Austria, Copyright (c) 2011-2017
--------------------------------------------------------------------------------
-- Description : 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- fixed_pkg resides in the library ieee since VHDL-2008 (QuestaSim backports
-- this to VHDL-93 too). However, Quartus (as of version 13.0sp1) still does
-- not have native support for ieee.fixed_pkg. Therefore, we provide the
-- VHDL-93 compatibility versions as part of this excercise. These must be
-- compiled into the are located in the library ieee_proposed. Include them in
-- your Config.tcl and don't forget to set the ExtraLibraries and TargetLibrary
-- parameters to compile them into the right library (ieee_proposed) with fhlow.
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
-- In future (when both QuestaSim and Quartus support the VHDL-2008
-- ieee.fixed_pkg) simply use:
--use ieee.fixed_float_types.all;
--use ieee.fixed_pkg.all;

use work.Global.all;

--------------------------------------------------------------------------------

entity tbDspFir is
end tbDspFir;

--------------------------------------------------------------------------------

architecture Bhv of tbDspFir is

  -- component generics
  constant cClkFrequency               : natural       := cDefaultClkFrequency;
  constant cIsLowPercentageOfDutyCycle : natural       := 65;
  constant cInResetDuration            : time          := 140 ns;
  constant cMclkFrequency              : natural       := 12E6;
  constant cSampleRate                 : natural       := cDefaultSampleRate;
  constant cAudioBitWidth              : natural       := cDefaultAudioBitWidth;
  constant cCoefWidth                  : natural       := 16;
  constant cB                          : aSetOfFactors := (-0.00013732910156250000,-0.00088119506835937500,0.00032806396484375000,0.00053405761718750000,-0.00053787231445312500,-0.00053405761718750000,0.00086975097656250000,0.00038909912109375000,-0.00119400024414063000,-0.00008392333984375000,0.00143814086914063000,-0.00035476684570312500,-0.00153350830078125000,0.00087356567382812500,0.00142669677734375000,-0.00138473510742188000,-0.00110244750976563000,0.00177764892578125000,0.00060653686523437500,-0.00197219848632813000,-0.00002670288085937500,0.00190353393554688000,-0.00051498413085937500,-0.00158691406250000000,0.00088119506835937500,0.00108718872070313000,-0.00097274780273437500,-0.00054168701171875000,0.00074005126953125000,0.00012207031250000000,-0.00022506713867187500,0.00001525878906250000,-0.00044631958007812500,0.00024414062500000000,0.00108337402343750000,-0.00091552734375000000,-0.00147247314453125000,0.00191879272460938000,0.00141906738281250000,-0.00305557250976563000,-0.00081253051757812500,0.00407409667968750000,-0.00032424926757812500,-0.00469970703125000000,0.00185012817382813000,0.00472259521484375000,-0.00349044799804688000,-0.00405120849609375000,0.00492477416992188000,0.00275039672851563000,-0.00583648681640625000,-0.00104522705078125000,0.00601196289062500000,-0.00071334838867187500,-0.00539779663085938000,0.00213623046875000000,0.00413131713867188000,-0.00288391113281250000,-0.00254440307617188000,0.00276565551757813000,0.00106430053710938000,-0.00179290771484375000,-0.00014495849609375000,0.00022506713867187500,0.00013351440429687500,0.00150299072265625000,-0.00116729736328125000,-0.00285720825195313000,0.00311660766601563000,0.00333786010742188000,-0.00559997558593750000,-0.00261306762695313000,0.00804138183593750000,0.00062942504882812500,-0.00980377197265625000,0.00234222412109375000,0.01034927368164060000,-0.00574874877929688000,-0.00940704345703125000,0.00886535644531250000,0.00704956054687500000,-0.01095581054687500000,-0.00373840332031250000,0.01148605346679690000,0.00024032592773437500,-0.01027297973632810000,0.00254440307617188000,0.00759887695312500000,-0.00377655029296875000,-0.00417327880859375000,0.00293350219726563000,0.00105667114257813000,0.00003051757812500000,0.00060653686523437500,-0.00457763671875000000,0.00017166137695312500,0.00964736938476563000,-0.00394821166992188000,-0.01381683349609380000,0.01063537597656250000,0.01557922363281250000,-0.01943588256835940000,-0.01369094848632810000,0.02891159057617190000,0.00746536254882813000,-0.03720855712890630000,0.00299453735351563000,0.04239654541015630000,-0.01672363281250000000,-0.04284286499023440000,0.03198623657226560000,0.03758621215820310000,-0.04655456542968750000,-0.02657318115234380000,0.05806732177734380000,0.01074600219726560000,-0.06448745727539060000,0.00806808471679688000,0.06446838378906250000,-0.02744293212890630000,-0.05765533447265630000,0.04475784301757810000,0.04475784301757810000,-0.05765533447265630000,-0.02744293212890630000,0.06446838378906250000,0.00806808471679688000,-0.06448745727539060000,0.01074600219726560000,0.05806732177734380000,-0.02657318115234380000,-0.04655456542968750000,0.03758621215820310000,0.03198623657226560000,-0.04284286499023440000,-0.01672363281250000000,0.04239654541015630000,0.00299453735351563000,-0.03720855712890630000,0.00746536254882813000,0.02891159057617190000,-0.01369094848632810000,-0.01943588256835940000,0.01557922363281250000,0.01063537597656250000,-0.01381683349609380000,-0.00394821166992188000,0.00964736938476563000,0.00017166137695312500,-0.00457763671875000000,0.00060653686523437500,0.00003051757812500000,0.00105667114257813000,0.00293350219726563000,-0.00417327880859375000,-0.00377655029296875000,0.00759887695312500000,0.00254440307617188000,-0.01027297973632810000,0.00024032592773437500,0.01148605346679690000,-0.00373840332031250000,-0.01095581054687500000,0.00704956054687500000,0.00886535644531250000,-0.00940704345703125000,-0.00574874877929688000,0.01034927368164060000,0.00234222412109375000,-0.00980377197265625000,0.00062942504882812500,0.00804138183593750000,-0.00261306762695313000,-0.00559997558593750000,0.00333786010742188000,0.00311660766601563000,-0.00285720825195313000,-0.00116729736328125000,0.00150299072265625000,0.00013351440429687500,0.00022506713867187500,-0.00014495849609375000,-0.00179290771484375000,0.00106430053710938000,0.00276565551757813000,-0.00254440307617188000,-0.00288391113281250000,0.00413131713867188000,0.00213623046875000000,-0.00539779663085938000,-0.00071334838867187500,0.00601196289062500000,-0.00104522705078125000,-0.00583648681640625000,0.00275039672851563000,0.00492477416992188000,-0.00405120849609375000,-0.00349044799804688000,0.00472259521484375000,0.00185012817382813000,-0.00469970703125000000,-0.00032424926757812500,0.00407409667968750000,-0.00081253051757812500,-0.00305557250976563000,0.00141906738281250000,0.00191879272460938000,-0.00147247314453125000,-0.00091552734375000000,0.00108337402343750000,0.00024414062500000000,-0.00044631958007812500,0.00001525878906250000,-0.00022506713867187500,0.00012207031250000000,0.00074005126953125000,-0.00054168701171875000,-0.00097274780273437500,0.00108718872070313000,0.00088119506835937500,-0.00158691406250000000,-0.00051498413085937500,0.00190353393554688000,-0.00002670288085937500,-0.00197219848632813000,0.00060653686523437500,0.00177764892578125000,-0.00110244750976563000,-0.00138473510742188000,0.00142669677734375000,0.00087356567382812500,-0.00153350830078125000,-0.00035476684570312500,0.00143814086914063000,-0.00008392333984375000,-0.00119400024414063000,0.00038909912109375000,0.00086975097656250000,-0.00053405761718750000,-0.00053787231445312500,0.00053405761718750000,0.00032806396484375000,-0.00088119506835937500,-0.00013732910156250000);
	--constant cB                          : aSetOfFactors := (0.25, 0.75, -0.25, 0.0, 0.125);
  --constant cB                          : aSetOfFactors := (-0.000152587890625, 0.00018310546875, 0.000152587890625, 0.000152587890625, 0.00018310546875, 0.000152587890625, 0.0001220703125, 0.00006103515625, 0.0, -0.000091552734375, -0.000213623046875, -0.00030517578125, -0.0003662109375, -0.0003662109375, -0.000335693359375, -0.000274658203125, -0.0001220703125, 0.00006103515625, 0.000244140625, 0.000457763671875, 0.0006103515625, 0.000732421875, 0.000732421875, 0.000640869140625, 0.000457763671875, 0.00018310546875, -0.000152587890625, -0.000518798828125, -0.0008544921875, -0.001129150390625, -0.001251220703125, -0.001251220703125, -0.00103759765625, -0.000701904296875, -0.000213623046875, 0.0003662109375, 0.000946044921875, 0.00146484375, 0.001861572265625, 0.00201416015625, 0.001922607421875, 0.001556396484375, 0.000946044921875, 0.000152587890625, -0.000732421875, -0.0015869140625, -0.0023193359375, -0.0028076171875, -0.002960205078125, -0.002716064453125, -0.002105712890625, -0.00115966796875, 0.0, 0.001251220703125, 0.00244140625, 0.00341796875, 0.00396728515625, 0.00408935546875, 0.003631591796875, 0.002685546875, 0.0013427734375, -0.00030517578125, -0.001983642578125, -0.0035400390625, -0.00469970703125, -0.005340576171875, -0.00531005859375, -0.00457763671875, -0.00323486328125, -0.001373291015625, 0.000762939453125, 0.0029296875, 0.004791259765625, 0.00616455078125, 0.00677490234375, 0.006561279296875, 0.0054931640625, 0.003631591796875, 0.001251220703125, -0.001434326171875, -0.0040283203125, -0.0062255859375, -0.0076904296875, -0.00823974609375, -0.00775146484375, -0.006256103515625, -0.003875732421875, -0.000946044921875, 0.00225830078125, 0.0052490234375, 0.007659912109375, 0.009185791015625, 0.00958251953125, 0.008758544921875, 0.006805419921875, 0.00390625, 0.00042724609375, -0.003204345703125, -0.006500244140625, -0.009063720703125, -0.010528564453125, -0.010711669921875, -0.009490966796875, -0.007080078125, -0.003692626953125, 0.000244140625, 0.004180908203125, 0.0076904296875, 0.010284423828125, 0.0115966796875, 0.011474609375, 0.0098876953125, 0.00701904296875, 0.00323486328125, -0.001007080078125, -0.005157470703125, -0.00872802734375, -0.011199951171875, -0.01226806640625, -0.011810302734375, -0.009857177734375, -0.00665283203125, -0.002593994140625, 0.0018310546875, 0.006011962890625, 0.00946044921875, 0.01171875, 0.01251220703125, 0.01171875, 0.00946044921875, 0.006011962890625, 0.0018310546875, -0.002593994140625, -0.00665283203125, -0.009857177734375, -0.011810302734375, -0.01226806640625, -0.011199951171875, -0.00872802734375, -0.005157470703125, -0.001007080078125, 0.00323486328125, 0.00701904296875, 0.0098876953125, 0.011474609375, 0.0115966796875, 0.010284423828125, 0.0076904296875, 0.004180908203125, 0.000244140625, -0.003692626953125, -0.007080078125, -0.009490966796875, -0.010711669921875, -0.010528564453125, -0.009063720703125, -0.006500244140625, -0.003204345703125, 0.00042724609375, 0.00390625, 0.006805419921875, 0.008758544921875, 0.00958251953125, 0.009185791015625, 0.007659912109375, 0.0052490234375, 0.00225830078125, -0.000946044921875, -0.003875732421875, -0.006256103515625, -0.00775146484375, -0.00823974609375, -0.0076904296875, -0.0062255859375, -0.0040283203125, -0.001434326171875, 0.001251220703125, 0.003631591796875, 0.0054931640625, 0.006561279296875, 0.00677490234375, 0.00616455078125, 0.004791259765625, 0.0029296875, 0.000762939453125, -0.001373291015625, -0.00323486328125, -0.00457763671875, -0.00531005859375, -0.005340576171875, -0.00469970703125, -0.0035400390625, -0.001983642578125, -0.00030517578125, 0.0013427734375, 0.002685546875, 0.003631591796875, 0.00408935546875, 0.00396728515625, 0.00341796875, 0.00244140625, 0.001251220703125, 0.0, -0.00115966796875, -0.002105712890625, -0.002716064453125, -0.002960205078125, -0.0028076171875, -0.0023193359375, -0.0015869140625, -0.000732421875, 0.000152587890625, 0.000946044921875, 0.001556396484375, 0.001922607421875, 0.00201416015625, 0.001861572265625, 0.00146484375, 0.000946044921875, 0.0003662109375, -0.000213623046875, -0.000701904296875, -0.00103759765625, -0.001251220703125, -0.001251220703125, -0.001129150390625, -0.0008544921875, -0.000518798828125, -0.000152587890625, 0.00018310546875, 0.000457763671875, 0.000640869140625, 0.000732421875, 0.000732421875, 0.0006103515625, 0.000457763671875, 0.000244140625, 0.00006103515625, -0.0001220703125, -0.000274658203125, -0.000335693359375, -0.0003662109375, -0.0003662109375, -0.00030517578125, -0.000213623046875, -0.000091552734375, 0.0, 0.00006103515625, 0.0001220703125, 0.000152587890625, 0.00018310546875, 0.000152587890625, 0.000152587890625, 0.00018310546875, -0.000152587890625);

  constant cWavName : string := "Wobble10Hz22050Hz100ms";

  constant cDryWavFileName    : string := "../../../../sounds/" & cWavName & ".wav";
  constant cWetWavFileName    : string := "Wet" & cWavName & ".wav";
  constant cWetRawWavFileName : string := "WetRawFile.raw";

  constant cRecordingDurationAftWaveEnd : time := 100 us;

  signal Clk                                : std_ulogic;
  signal nResetAsync                        : std_ulogic;
  signal DdryL, DdryR, DwetL, DwetR         : aAudioData(0 downto -(cAudioBitWidth-1));
  signal ValDryL, ValDryR, ValWetL, ValWetR : std_ulogic;
  signal WaveAtEnd                          : boolean := false;
  signal ADClrc                             : std_ulogic;
  signal Mclk                               : std_ulogic;
  signal Bclk                               : std_ulogic;

begin

  TheWavToPar : entity work.WavToPar
    generic map (
      gWaveFileName  => cDryWavFileName,
      gSampleRate    => cSampleRate,
      gAudioBitWidth => cAudioBitWidth)
    port map (
      iClk       => Clk,
      oDL        => DdryL,
      oDR        => DdryR,
      oValL      => ValDryL,
      oValR      => ValDryR,
      oWaveAtEnd => WaveAtEnd,
      iLrc       => ADClrc);

  FirInstance : entity work.DspFir(RtlRam)
    generic map (
      gAudioBitWidth => cAudioBitWidth,
      gCoefWidth     => cCoefWidth,
      gB             => cB
      )
    port map (
      iClk         => Clk,
      inResetAsync => nResetAsync,
      iDdry        => DdryL,
      iValDry      => ValDryL,
      oDwet        => DwetL,
      oValWet      => ValWetL);

  DwetR   <= DdryR;
  ValWetR <= ValDryR;

  TheParToWav : entity work.ParToWav
    generic map (
      gWavFileName                 => cWetWavFileName,
      gRawWavFileName              => cWetRawWavFileName,
      gRecordingDurationAftWaveEnd => cRecordingDurationAftWaveEnd,
      gFormatTag                   => open,
      gAudioBitWidth               => open,
      gChannels                    => open,
      gSampleRate                  => cDefaultSampleRate)
    port map (
      iClk       => Clk,
      iDL        => DwetL,
      iDR        => DwetR,
      iValL      => ValWetL,
      iValR      => ValWetR,
      iWaveAtEnd => WaveAtEnd);

  GenClks : entity work.ClkMaster
    generic map (
      gClkFrequency  => cClkFrequency,
      gMclkFrequency => cMclkFrequency,
      gSampleRate    => cSampleRate)
    port map (
      iClk         => Clk,
      inResetAsync => nResetAsync,
      oMclk        => Mclk,
      oBclk        => Bclk,
      oADClrc      => ADClrc);

  ClkGen : entity work.Oscillator
    generic map (
      gFrequency                  => cClkFrequency,
      gIsLowPercentageOfDutyCycle => cIsLowPercentageOfDutyCycle)
    port map (
      oRectangleWave => Clk);

  -- reset generation
  PwrOnResetSource : entity work.PwrOnReset
    generic map (
      gInResetDuration => cInResetDuration,
      gResetLevel      => cResetActive)
    port map (
      onResetAsync => nResetAsync);

end Bhv;
